`default_nettype none

// `define SIN
